LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY   IS
  GENERIC();
  PORT();
END ;

ARCHITECTURE arch OF  IS

  BEGIN

  
END arch;
